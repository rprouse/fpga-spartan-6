
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity BlinkLeds_HDL is
    Port ( CLOCK_IN : in  STD_LOGIC;
           RESET : in  STD_LOGIC;
           OUT_HIGH : out  STD_LOGIC;
           OUT_LOW : out  STD_LOGIC);
end BlinkLeds_HDL;

architecture Behavioral of BlinkLeds_HDL is

begin


end Behavioral;

